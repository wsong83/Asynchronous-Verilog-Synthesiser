module test_module;
   wire o;
   assign o = 3;
   
endmodule // test

