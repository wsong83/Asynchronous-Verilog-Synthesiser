module test_module (o);
   output [2:0] o;
   wire [2:0]   o;
   reg [4+25:4'd35] sig, tmp;
   
   assign o = {3'b11};
   
endmodule // test

module test_module;
endmodule // test_module

/*
 
 

