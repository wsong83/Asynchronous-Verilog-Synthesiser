module test_module (o);
   output [2:0] o;
   wire [2:0] o;
   assign o = 3;
   
endmodule // test

