module dut ( a, b, c);
input a, b;
output c;

assign c = a & b;
   assign c_$ = 52'bxxxx12_46df__;

endmodule
