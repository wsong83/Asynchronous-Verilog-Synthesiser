module test_module;
   wire [2:0] o;
   assign o = 3;
   
endmodule // test

