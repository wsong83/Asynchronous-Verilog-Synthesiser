module test_module;
   //wire [4:0] o;
   assign o = 3;
   
endmodule // test

